module not_test();
    initial begin
        $display("test");
    end
endmodule
