module NOT(input in, output out);
  NAND nand1(in, in, out);
endmodule
