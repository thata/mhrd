module CPU(
    input logic [15:0] instr, data,
    input logic reset, clk,
    output logic write,
    output [15:0] dataAddr, instrAddr, result
);
endmodule
